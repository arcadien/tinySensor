.title KiCad schematic
R2 +3V3 /SDA 4,7k
R3 +3V3 /SCL 4,7k
U1 +3V3 NC_01 /LED_OUT NC_02 NC_03 /TX_RADIO /SDA NC_04 /SCL NC_05 NC_06 NC_07 NC_08 GND ATtiny84A-PU
R1 GND Net-_D1-Pad1_ 1k
D1 Net-_D1-Pad1_ /LED_OUT LED
J1 +3V3 GND /TX_RADIO RADIO
J3 +3V3 GND /SCL /SDA NC_09 GND NC_10 BMP/BME breakout
J2 +BATT GND +3V3 NC_11 DCDC converter
C1 +3V3 GND 10u
C2 GND +3V3 100n
.end
